module mult (
	input [15:0] a, b, 
	output [15:0] product 

);

assign product = a * b;

endmodule 
